//=============================================================================
// Module Name: sdcard_data_engine
//=============================================================================
// Description: SD Data Engine for SD Card Controller
//              Handles data block transmission/reception with CRC checking
//              and FIFO management for high-performance data transfer
//
// Features:
// - Data block transmission and reception
// - CRC16 generation and checking for data
// - FIFO management and flow control
// - Multiple data width support (1, 4, 8 bits)
// - Performance optimization
// - Error detection and recovery
// - DMA interface support
//
// Author: Vyges Development Team
// License: Apache-2.0
//=============================================================================

module sdcard_data_engine #(
    parameter int SDCARD_DATA_WIDTH = 4,
    parameter int FIFO_DEPTH = 512
) (
    // Clock and Reset
    input  logic                    PCLK_i,           // APB clock
    input  logic                    PRESETn_i,        // APB reset, active low
    
    // SD Card Interface
    input  logic                   sd_clk_o,          // SD card clock
    inout  logic [SDCARD_DATA_WIDTH-1:0] sd_dat_io,       // SD data lines
    
    // Data Interface
    input  logic [31:0]            data_in,           // Data input
    output logic [31:0]            data_out,          // Data output
    input  logic                   data_valid,        // Data valid
    output logic                   data_ready,        // Data ready
    input  logic                   data_start,        // Data start
    output logic                   data_busy,         // Data busy
    output logic                   data_done,         // Data done
    output logic [15:0]            data_crc,          // Data CRC
    output logic                   data_crc_error,    // Data CRC error
    
    // FIFO Interface
    input  logic [31:0]            fifo_data_in,      // FIFO data input
    output logic [31:0]            fifo_data_out,     // FIFO data output
    input  logic                   fifo_write,        // FIFO write enable
    output logic                   fifo_read,         // FIFO read enable
    input  logic                   fifo_full,         // FIFO full
    input  logic                   fifo_empty,        // FIFO empty
    input  logic [9:0]             fifo_count,        // FIFO count
    
    // Clock Interface
    input  logic                   clk_enable,        // Clock enable
    input  logic [15:0]            clk_divider,       // Clock divider
    
    // Power and Security Interface
    input  logic [1:0]             power_state,       // Power state
    input  logic                   security_lock,     // Security lock
    input  logic                   access_granted,    // Access granted
    
    // Error Interface
    input  logic [15:0]            error_status,      // Error status
    output logic                   error_clear        // Error clear
);

    // Data engine state machine states
    typedef enum logic [3:0] {
        DATA_IDLE = 4'b0000,
        DATA_SETUP = 4'b0001,
        DATA_TX_START = 4'b0010,
        DATA_TX_BLOCK = 4'b0011,
        DATA_TX_CRC = 4'b0100,
        DATA_TX_END = 4'b0101,
        DATA_RX_START = 4'b0110,
        DATA_RX_BLOCK = 4'b0111,
        DATA_RX_CRC = 4'b1000,
        DATA_RX_END = 4'b1001,
        DATA_COMPLETE = 4'b1010,
        DATA_ERROR = 4'b1011,
        DATA_TIMEOUT = 4'b1100
    } data_state_t;
    
    data_state_t data_state, data_next_state;
    
    // Internal signals
    logic [31:0]                   tx_data;           // Transmit data
    logic [31:0]                   rx_data;           // Receive data
    logic [15:0]                   tx_crc;            // Transmit CRC
    logic [15:0]                   rx_crc;            // Receive CRC
    logic [15:0]                   calc_crc;          // Calculated CRC
    logic [9:0]                    byte_counter;      // Byte counter
    logic [7:0]                    bit_counter;       // Bit counter
    logic [15:0]                   timeout_counter;   // Timeout counter
    logic [15:0]                   timeout_limit;     // Timeout limit
    logic [SDCARD_DATA_WIDTH-1:0]      data_out_bits;     // Data output bits
    logic [SDCARD_DATA_WIDTH-1:0]      data_in_bits;      // Data input bits
    logic                          data_out_en;       // Data output enable
    logic                          crc_valid;         // CRC valid
    logic                          timeout_expired;   // Timeout expired
    logic                          is_write;          // Write operation
    logic                          is_read;           // Read operation
    logic [11:0]                   block_size;        // Block size in bytes
    
    // Data width configuration
    localparam [1:0] DATA_WIDTH_1BIT = 2'b00;
    localparam [1:0] DATA_WIDTH_4BIT = 2'b01;
    localparam [1:0] DATA_WIDTH_8BIT = 2'b10;
    
    // Data state machine
    always_ff @(posedge PCLK_i or negedge PRESETn_i) begin
        if (!PRESETn_i) begin
            data_state <= DATA_IDLE;
        end else begin
            data_state <= data_next_state;
        end
    end
    
    // Data state machine next state logic
    always_comb begin
        data_next_state = data_state;
        
        case (data_state)
            DATA_IDLE: begin
                if (data_start && clk_enable && !security_lock && access_granted) begin
                    if (data_valid) begin
                        data_next_state = DATA_TX_START;
                    end else begin
                        data_next_state = DATA_RX_START;
                    end
                end
            end
            
            DATA_SETUP: begin
                data_next_state = is_write ? DATA_TX_START : DATA_RX_START;
            end
            
            DATA_TX_START: begin
                data_next_state = DATA_TX_BLOCK;
            end
            
            DATA_TX_BLOCK: begin
                if (byte_counter >= block_size) begin
                    data_next_state = DATA_TX_CRC;
                end
            end
            
            DATA_TX_CRC: begin
                if (bit_counter == 8'd15) begin
                    data_next_state = DATA_TX_END;
                end
            end
            
            DATA_TX_END: begin
                data_next_state = DATA_COMPLETE;
            end
            
            DATA_RX_START: begin
                if (timeout_expired) begin
                    data_next_state = DATA_TIMEOUT;
                end else if (data_in_bits != 4'hF) begin
                    data_next_state = DATA_RX_BLOCK;
                end
            end
            
            DATA_RX_BLOCK: begin
                if (byte_counter >= block_size) begin
                    data_next_state = DATA_RX_CRC;
                end
            end
            
            DATA_RX_CRC: begin
                if (bit_counter == 8'd15) begin
                    data_next_state = DATA_RX_END;
                end
            end
            
            DATA_RX_END: begin
                if (crc_valid) begin
                    data_next_state = DATA_COMPLETE;
                else begin
                    data_next_state = DATA_ERROR;
                end
            end
            
            DATA_COMPLETE: begin
                data_next_state = DATA_IDLE;
            end
            
            DATA_ERROR: begin
                data_next_state = DATA_IDLE;
            end
            
            DATA_TIMEOUT: begin
                data_next_state = DATA_IDLE;
            end
            
            default: begin
                data_next_state = DATA_IDLE;
            end
        endcase
    end
    
    // CRC16 calculation for data
    function automatic [15:0] calc_crc16;
        input [7:0] data;
        input [15:0] crc_in;
        reg [15:0] crc;
        integer i;
        begin
            crc = crc_in;
            for (i = 7; i >= 0; i = i - 1) begin
                crc = {crc[14:0], 1'b0} ^ (crc[15] ^ data[i] ? 16'h1021 : 16'h0000);
            end
            calc_crc16 = crc;
        end
    endfunction
    
    // Data control logic
    always_ff @(posedge PCLK_i or negedge PRESETn_i) begin
        if (!PRESETn_i) begin
            data_busy <= 1'b0;
            data_done <= 1'b0;
            data_crc_error <= 1'b0;
            data_ready <= 1'b1;
            data_out <= 32'h0;
            data_crc <= 16'h0;
            tx_data <= 32'h0;
            rx_data <= 32'h0;
            tx_crc <= 16'h0;
            rx_crc <= 16'h0;
            byte_counter <= 10'h0;
            bit_counter <= 8'h0;
            timeout_counter <= 16'h0;
            timeout_limit <= 16'hFFFF;
            data_out_bits <= {SDCARD_DATA_WIDTH{1'b1}};
            data_out_en <= 1'b0;
            crc_valid <= 1'b0;
            timeout_expired <= 1'b0;
            is_write <= 1'b0;
            is_read <= 1'b0;
            block_size <= 12'h200; // 512 bytes default
            error_clear <= 1'b0;
            fifo_read <= 1'b0;
        end else begin
            // Default values
            data_done <= 1'b0;
            data_crc_error <= 1'b0;
            error_clear <= 1'b0;
            fifo_read <= 1'b0;
            
            case (data_state)
                DATA_IDLE: begin
                    data_busy <= 1'b0;
                    data_ready <= 1'b1;
                    data_out_en <= 1'b0;
                    byte_counter <= 10'h0;
                    bit_counter <= 8'h0;
                    timeout_counter <= 16'h0;
                    timeout_expired <= 1'b0;
                    crc_valid <= 1'b0;
                    tx_crc <= 16'h0;
                    rx_crc <= 16'h0;
                    
                    if (data_start) begin
                        is_write <= data_valid;
                        is_read <= !data_valid;
                        block_size <= 12'h200; // Default 512 bytes
                        timeout_limit <= 16'hFFFF;
                    end
                end
                
                DATA_SETUP: begin
                    data_busy <= 1'b1;
                    data_ready <= 1'b0;
                end
                
                DATA_TX_START: begin
                    if (is_write) begin
                        tx_data <= data_in;
                        data_out_en <= 1'b1;
                    end
                end
                
                DATA_TX_BLOCK: begin
                    // Transmit data bytes
                    if (byte_counter < block_size) begin
                        case (SDCARD_DATA_WIDTH)
                            1: begin
                                data_out_bits[0] <= tx_data[31 - byte_counter];
                            end
                            4: begin
                                data_out_bits <= tx_data[31 - byte_counter*4 -: 4];
                            end
                            8: begin
                                data_out_bits <= tx_data[31 - byte_counter*8 -: 8];
                            end
                            default: begin
                                data_out_bits <= tx_data[31 - byte_counter*4 -: 4];
                            end
                        endcase
                        
                        // Update CRC
                        tx_crc <= calc_crc16(tx_data[31 - byte_counter*8 -: 8], tx_crc);
                        byte_counter <= byte_counter + 10'h1;
                    end
                end
                
                DATA_TX_CRC: begin
                    // Transmit CRC
                    data_out_bits <= tx_crc[15 - bit_counter];
                    bit_counter <= bit_counter + 8'h1;
                end
                
                DATA_TX_END: begin
                    data_out_en <= 1'b0;
                    data_crc <= tx_crc;
                end
                
                DATA_RX_START: begin
                    data_out_en <= 1'b0;
                    timeout_counter <= timeout_counter + 16'h1;
                    timeout_expired <= (timeout_counter >= timeout_limit);
                end
                
                DATA_RX_BLOCK: begin
                    // Receive data bytes
                    if (byte_counter < block_size) begin
                        case (SDCARD_DATA_WIDTH)
                            1: begin
                                rx_data[31 - byte_counter] <= data_in_bits[0];
                            end
                            4: begin
                                rx_data[31 - byte_counter*4 -: 4] <= data_in_bits;
                            end
                            8: begin
                                rx_data[31 - byte_counter*8 -: 8] <= data_in_bits;
                            end
                            default: begin
                                rx_data[31 - byte_counter*4 -: 4] <= data_in_bits;
                            end
                        endcase
                        
                        // Update CRC
                        rx_crc <= calc_crc16(rx_data[31 - byte_counter*8 -: 8], rx_crc);
                        byte_counter <= byte_counter + 10'h1;
                    end
                end
                
                DATA_RX_CRC: begin
                    // Receive CRC
                    rx_crc[15 - bit_counter] <= data_in_bits[0];
                    bit_counter <= bit_counter + 8'h1;
                end
                
                DATA_RX_END: begin
                    // Check CRC
                    calc_crc <= calc_crc16(rx_data[31 - byte_counter*8 -: 8], rx_crc);
                    crc_valid <= (calc_crc16(rx_data[31 - byte_counter*8 -: 8], rx_crc) == rx_crc);
                end
                
                DATA_COMPLETE: begin
                    data_done <= 1'b1;
                    data_busy <= 1'b0;
                    data_ready <= 1'b1;
                    
                    if (is_read) begin
                        data_out <= rx_data;
                        data_crc <= rx_crc;
                    end
                end
                
                DATA_ERROR: begin
                    data_crc_error <= 1'b1;
                    data_busy <= 1'b0;
                    data_ready <= 1'b1;
                    error_clear <= 1'b1;
                end
                
                DATA_TIMEOUT: begin
                    data_busy <= 1'b0;
                    data_ready <= 1'b1;
                    error_clear <= 1'b1;
                end
                
                default: begin
                    // No action
                end
            endcase
        end
    end
    
    // SD data lines control
    genvar i;
    generate
        for (i = 0; i < SDCARD_DATA_WIDTH; i = i + 1) begin : data_lines
            assign sd_dat_io[i] = data_out_en ? data_out_bits[i] : 1'bz;
            assign data_in_bits[i] = sd_dat_io[i];
        end
    endgenerate
    
    // FIFO interface
    always_ff @(posedge PCLK_i) begin
        if (fifo_write && !fifo_full) begin
            // Write data to FIFO
        end
        
        if (fifo_read && !fifo_empty) begin
            // Read data from FIFO
            fifo_data_out <= fifo_data_in;
        end
    end
    
    // Assertions for data protocol compliance
    // synthesis translate_off
    property data_start_condition;
        @(posedge PCLK_i) data_start |-> ##1 data_busy;
    endproperty
    
    property data_completion;
        @(posedge PCLK_i) data_busy |-> ##[1:10000] (data_done || data_crc_error);
    endproperty
    
    property data_crc_error_valid;
        @(posedge PCLK_i) data_crc_error |-> !data_done;
    endproperty
    
    property fifo_overflow_protection;
        @(posedge PCLK_i) fifo_full |-> !fifo_write;
    endproperty
    
    property fifo_underflow_protection;
        @(posedge PCLK_i) fifo_empty |-> !fifo_read;
    endproperty
    
    data_start_condition_check: assert property (data_start_condition)
        else $error("Data start condition violation");
    
    data_completion_check: assert property (data_completion)
        else $error("Data completion violation");
    
    data_crc_error_valid_check: assert property (data_crc_error_valid)
        else $error("Data CRC error validity violation");
    
    fifo_overflow_protection_check: assert property (fifo_overflow_protection)
        else $error("FIFO overflow protection violation");
    
    fifo_underflow_protection_check: assert property (fifo_underflow_protection)
        else $error("FIFO underflow protection violation");
    // synthesis translate_on

endmodule 