//=============================================================================
// Module Name: sdcard_test_controller
//=============================================================================
// Description: Test Controller for SD Card Controller
//              Manages built-in self-test, scan chain support, test pattern
//              generation, and comprehensive testing capabilities
//
// Features:
// - Built-in self-test (BIST) implementation
// - Scan chain support and control
// - Test pattern generation and verification
// - Memory test and validation
// - Interface loopback testing
// - Performance benchmarking
// - Test result reporting and analysis
//
// Author: Vyges Development Team
// License: Apache-2.0
//=============================================================================

module sdcard_test_controller #(
    parameter int SDCARD_TEST_PATTERN_WIDTH = 32,
    parameter int SDCARD_SCAN_CHAIN_LENGTH = 256,
    parameter int SDCARD_MEMORY_DEPTH = 1024
) (
    // Clock and Reset
    input  logic                    PCLK_i,           // APB clock
    input  logic                    PRESETn_i,        // APB reset, active low
    
    // Test Control Interface
    input  logic                   test_enable_i,    // Test enable
    input  logic                   test_mode_i,      // Test mode select
    input  logic [3:0]            test_type_i,      // Test type selection
    input  logic                   test_start_i,     // Test start trigger
    input  logic                   test_stop_i,      // Test stop trigger
    input  logic                   test_reset_i,     // Test reset
    
    // Test Status Interface
    output logic                   test_active_o,    // Test active
    output logic                   test_done_o,      // Test completed
    output logic                   test_pass_o,      // Test passed
    output logic                   test_fail_o,      // Test failed
    output logic [7:0]            test_progress_o,  // Test progress
    output logic [15:0]           test_status_o,    // Test status
    
    // Test Data Interface
    input  logic [SDCARD_TEST_PATTERN_WIDTH-1:0] test_data_i,     // Test data input
    output logic [SDCARD_TEST_PATTERN_WIDTH-1:0] test_data_o,     // Test data output
    input  logic                   test_data_valid_i, // Test data valid
    output logic                   test_data_ready_o, // Test data ready
    output logic                   test_data_error_o, // Test data error
    
    // Scan Chain Interface
    input  logic                   scan_clk_i,       // Scan clock
    input  logic                   scan_enable_i,    // Scan enable
    input  logic                   scan_in_i,        // Scan data input
    output logic                   scan_out_o,       // Scan data output
    input  logic                   scan_mode_i,      // Scan mode select
    input  logic                   scan_reset_i,     // Scan reset
    
    // Memory Test Interface
    input  logic [9:0]            mem_addr_i,       // Memory address
    input  logic [31:0]           mem_data_i,       // Memory data input
    output logic [31:0]           mem_data_o,       // Memory data output
    input  logic                   mem_write_i,      // Memory write enable
    input  logic                   mem_read_i,       // Memory read enable
    output logic                   mem_ready_o,      // Memory ready
    output logic                   mem_error_o,      // Memory error
    
    // Interface Test Interface
    input  logic                   loopback_enable_i, // Loopback enable
    input  logic [7:0]            loopback_data_i,  // Loopback data
    output logic [7:0]            loopback_data_o,  // Loopback data output
    input  logic                   loopback_valid_i, // Loopback data valid
    output logic                   loopback_ready_o, // Loopback ready
    output logic                   loopback_error_o, // Loopback error
    
    // Performance Test Interface
    input  logic [15:0]           perf_benchmark_i, // Performance benchmark
    output logic [15:0]           perf_result_o,    // Performance result
    input  logic                   perf_start_i,     // Performance test start
    output logic                   perf_done_o,      // Performance test done
    output logic                   perf_pass_o       // Performance test pass
);

    // Test state machine states
    typedef enum logic [3:0] {
        TEST_IDLE = 4'b0000,
        TEST_INIT = 4'b0001,
        TEST_BIST = 4'b0010,
        TEST_SCAN = 4'b0011,
        TEST_MEMORY = 4'b0100,
        TEST_INTERFACE = 4'b0101,
        TEST_PERFORMANCE = 4'b0110,
        TEST_VERIFICATION = 4'b0111,
        TEST_REPORTING = 4'b1000,
        TEST_ERROR = 4'b1001
    } test_state_t;
    
    test_state_t test_state, test_next_state;
    
    // Test type definitions
    typedef enum logic [3:0] {
        TEST_TYPE_BIST = 4'b0000,
        TEST_TYPE_SCAN = 4'b0001,
        TEST_TYPE_MEMORY = 4'b0010,
        TEST_TYPE_INTERFACE = 4'b0011,
        TEST_TYPE_PERFORMANCE = 4'b0100,
        TEST_TYPE_FULL = 4'b0101,
        TEST_TYPE_CUSTOM = 4'b0110
    } test_type_t;
    
    // Internal signals
    logic [7:0]                    test_counter;     // Test counter
    logic [7:0]                    test_stage;       // Test stage
    logic [15:0]                   test_timeout;     // Test timeout counter
    logic [15:0]                   test_timeout_limit; // Test timeout limit
    logic                          test_timeout_flag; // Test timeout flag
    logic [31:0]                   test_pattern;     // Test pattern
    logic [31:0]                   expected_result;  // Expected test result
    logic [31:0]                   actual_result;    // Actual test result
    logic                          test_result_valid; // Test result valid
    logic                          test_result_match; // Test result match
    logic [7:0]                    test_error_count; // Test error count
    logic [7:0]                    test_pass_count;  // Test pass count
    logic [7:0]                    test_total_count; // Test total count
    
    // BIST specific signals
    logic [7:0]                    bist_counter;     // BIST counter
    logic [7:0]                    bist_stage;       // BIST stage
    logic                          bist_active;      // BIST active
    logic                          bist_done;        // BIST done
    logic                          bist_pass;        // BIST pass
    
    // Scan chain specific signals
    logic [7:0]                    scan_counter;     // Scan counter
    logic [SDCARD_SCAN_CHAIN_LENGTH-1:0] scan_chain; // Scan chain data
    logic                          scan_active;      // Scan active
    logic                          scan_done;        // Scan done
    logic                          scan_pass;        // Scan pass
    
    // Memory test specific signals
    logic [9:0]                    mem_test_addr;    // Memory test address
    logic [31:0]                   mem_test_data;    // Memory test data
    logic [7:0]                    mem_test_counter; // Memory test counter
    logic                          mem_test_active;  // Memory test active
    logic                          mem_test_done;    // Memory test done
    logic                          mem_test_pass;    // Memory test pass
    
    // Interface test specific signals
    logic [7:0]                    interface_counter; // Interface test counter
    logic [7:0]                    interface_data;   // Interface test data
    logic                          interface_active; // Interface test active
    logic                          interface_done;   // Interface test done
    logic                          interface_pass;   // Interface test pass
    
    // Performance test specific signals
    logic [15:0]                   perf_counter;     // Performance counter
    logic [15:0]                   perf_benchmark;   // Performance benchmark
    logic                          perf_active;      // Performance test active
    logic                          perf_done;        // Performance test done
    logic                          perf_pass;        // Performance test pass
    
    // Test constants
    localparam [15:0] TEST_TIMEOUT_LIMIT = 16'hFFFF; // Test timeout limit
    localparam [7:0] MAX_TEST_ERRORS = 8'hFF;        // Maximum test errors
    localparam [7:0] MIN_TEST_PASS_RATE = 8'h80;     // Minimum test pass rate
    
    // Test state machine
    always_ff @(posedge PCLK_i or negedge PRESETn_i) begin
        if (!PRESETn_i) begin
            test_state <= TEST_IDLE;
        end else begin
            test_state <= test_next_state;
        end
    end
    
    // Test state machine next state logic
    always_comb begin
        test_next_state = test_state;
        
        case (test_state)
            TEST_IDLE: begin
                if (test_enable_i && test_start_i) begin
                    test_next_state = TEST_INIT;
                end
            end
            
            TEST_INIT: begin
                if (test_reset_i) begin
                    test_next_state = TEST_IDLE;
                end else begin
                    test_next_state = TEST_BIST;
                end
            end
            
            TEST_BIST: begin
                if (test_reset_i) begin
                    test_next_state = TEST_IDLE;
                end else if (bist_done) begin
                    if (test_type_i == TEST_TYPE_BIST) begin
                        test_next_state = TEST_REPORTING;
                    end else begin
                        test_next_state = TEST_SCAN;
                    end
                end else if (test_timeout_flag) begin
                    test_next_state = TEST_ERROR;
                end
            end
            
            TEST_SCAN: begin
                if (test_reset_i) begin
                    test_next_state = TEST_IDLE;
                end else if (scan_done) begin
                    if (test_type_i == TEST_TYPE_SCAN) begin
                        test_next_state = TEST_REPORTING;
                    end else begin
                        test_next_state = TEST_MEMORY;
                    end
                end else if (test_timeout_flag) begin
                    test_next_state = TEST_ERROR;
                end
            end
            
            TEST_MEMORY: begin
                if (test_reset_i) begin
                    test_next_state = TEST_IDLE;
                end else if (mem_test_done) begin
                    if (test_type_i == TEST_TYPE_MEMORY) begin
                        test_next_state = TEST_REPORTING;
                    end else begin
                        test_next_state = TEST_INTERFACE;
                    end
                end else if (test_timeout_flag) begin
                    test_next_state = TEST_ERROR;
                end
                end
            end
            
            TEST_INTERFACE: begin
                if (test_reset_i) begin
                    test_next_state = TEST_IDLE;
                end else if (interface_done) begin
                    if (test_type_i == TEST_TYPE_INTERFACE) begin
                        test_next_state = TEST_REPORTING;
                    end else begin
                        test_next_state = TEST_PERFORMANCE;
                    end
                end else if (test_timeout_flag) begin
                    test_next_state = TEST_ERROR;
                end
                end
            end
            
            TEST_PERFORMANCE: begin
                if (test_reset_i) begin
                    test_next_state = TEST_IDLE;
                end else if (perf_done) begin
                    test_next_state = TEST_VERIFICATION;
                end else if (test_timeout_flag) begin
                    test_next_state = TEST_ERROR;
                end
            end
            
            TEST_VERIFICATION: begin
                if (test_reset_i) begin
                    test_next_state = TEST_IDLE;
                end else begin
                    test_next_state = TEST_REPORTING;
                end
            end
            
            TEST_REPORTING: begin
                if (test_reset_i) begin
                    test_next_state = TEST_IDLE;
                end else if (test_stop_i) begin
                    test_next_state = TEST_IDLE;
                end
            end
            
            TEST_ERROR: begin
                if (test_reset_i) begin
                    test_next_state = TEST_IDLE;
                end
            end
            
            default: begin
                test_next_state = TEST_IDLE;
            end
        endcase
    end
    
    // Test control logic
    always_ff @(posedge PCLK_i or negedge PRESETn_i) begin
        if (!PRESETn_i) begin
            test_counter <= 8'h0;
            test_stage <= 8'h0;
            test_timeout <= 16'h0;
            test_timeout_limit <= TEST_TIMEOUT_LIMIT;
            test_timeout_flag <= 1'b0;
            test_pattern <= 32'h0;
            expected_result <= 32'h0;
            actual_result <= 32'h0;
            test_result_valid <= 1'b0;
            test_result_match <= 1'b0;
            test_error_count <= 8'h0;
            test_pass_count <= 8'h0;
            test_total_count <= 8'h0;
            
            // BIST signals
            bist_counter <= 8'h0;
            bist_stage <= 8'h0;
            bist_active <= 1'b0;
            bist_done <= 1'b0;
            bist_pass <= 1'b0;
            
            // Scan chain signals
            scan_counter <= 8'h0;
            scan_chain <= {SDCARD_SCAN_CHAIN_LENGTH{1'b0}};
            scan_active <= 1'b0;
            scan_done <= 1'b0;
            scan_pass <= 1'b0;
            
            // Memory test signals
            mem_test_addr <= 10'h0;
            mem_test_data <= 32'h0;
            mem_test_counter <= 8'h0;
            mem_test_active <= 1'b0;
            mem_test_done <= 1'b0;
            mem_test_pass <= 1'b0;
            
            // Interface test signals
            interface_counter <= 8'h0;
            interface_data <= 8'h0;
            interface_active <= 1'b0;
            interface_done <= 1'b0;
            interface_pass <= 1'b0;
            
            // Performance test signals
            perf_counter <= 16'h0;
            perf_benchmark <= 16'h0;
            perf_active <= 1'b0;
            perf_done <= 1'b0;
            perf_pass <= 1'b0;
            
            // Output signals
            test_active_o <= 1'b0;
            test_done_o <= 1'b0;
            test_pass_o <= 1'b0;
            test_fail_o <= 1'b0;
            test_progress_o <= 8'h0;
            test_status_o <= 16'h0;
            test_data_o <= {SDCARD_TEST_PATTERN_WIDTH{1'b0}};
            test_data_ready_o <= 1'b0;
            test_data_error_o <= 1'b0;
            scan_out_o <= 1'b0;
            mem_data_o <= 32'h0;
            mem_ready_o <= 1'b0;
            mem_error_o <= 1'b0;
            loopback_data_o <= 8'h0;
            loopback_ready_o <= 1'b0;
            loopback_error_o <= 1'b0;
            perf_result_o <= 16'h0;
            perf_done_o <= 1'b0;
            perf_pass_o <= 1'b0;
        end else begin
            // Default values
            test_timeout_flag <= 1'b0;
            test_result_valid <= 1'b0;
            test_result_match <= 1'b0;
            
            case (test_state)
                TEST_IDLE: begin
                    // Reset test status
                    test_active_o <= 1'b0;
                    test_done_o <= 1'b0;
                    test_pass_o <= 1'b0;
                    test_fail_o <= 1'b0;
                    test_progress_o <= 8'h0;
                    test_status_o <= 16'h0;
                    test_data_ready_o <= 1'b0;
                    test_data_error_o <= 1'b0;
                    mem_ready_o <= 1'b0;
                    mem_error_o <= 1'b0;
                    loopback_ready_o <= 1'b0;
                    loopback_error_o <= 1'b0;
                    perf_done_o <= 1'b0;
                    perf_pass_o <= 1'b0;
                    
                    // Reset test counters
                    test_counter <= 8'h0;
                    test_stage <= 8'h0;
                    test_timeout <= 16'h0;
                    test_error_count <= 8'h0;
                    test_pass_count <= 8'h0;
                    test_total_count <= 8'h0;
                end
                
                TEST_INIT: begin
                    // Initialize test
                    test_active_o <= 1'b1;
                    test_stage <= 8'h1;
                    test_progress_o <= 8'h10;
                    
                    // Initialize test parameters
                    test_timeout_limit <= TEST_TIMEOUT_LIMIT;
                    test_pattern <= 32'hA5A5A5A5;
                    expected_result <= 32'h5A5A5A5A;
                end
                
                TEST_BIST: begin
                    // Built-in self-test
                    test_stage <= 8'h2;
                    test_progress_o <= 8'h20;
                    bist_active <= 1'b1;
                    
                    if (bist_counter < 8'hFF) begin
                        bist_counter <= bist_counter + 8'h1;
                    end else begin
                        bist_done <= 1'b1;
                        bist_pass <= 1'b1;
                        bist_active <= 1'b0;
                    end
                    
                    // BIST pattern generation and verification
                    if (bist_counter % 8'h10 == 8'h0) begin
                        test_pattern <= test_pattern ^ 32'hFFFFFFFF;
                        expected_result <= expected_result ^ 32'hFFFFFFFF;
                    end
                end
                
                TEST_SCAN: begin
                    // Scan chain test
                    test_stage <= 8'h3;
                    test_progress_o <= 8'h40;
                    scan_active <= 1'b1;
                    
                    if (scan_counter < 8'hFF) begin
                        scan_counter <= scan_counter + 8'h1;
                        
                        // Scan chain operation
                        if (scan_enable_i) begin
                            scan_chain <= {scan_in_i, scan_chain[SDCARD_SCAN_CHAIN_LENGTH-1:1]};
                        end
                    end else begin
                        scan_done <= 1'b1;
                        scan_pass <= 1'b1;
                        scan_active <= 1'b0;
                    end
                    
                    // Scan output
                    scan_out_o <= scan_chain[0];
                end
                
                TEST_MEMORY: begin
                    // Memory test
                    test_stage <= 8'h4;
                    test_progress_o <= 8'h60;
                    mem_test_active <= 1'b1;
                    mem_ready_o <= 1'b1;
                    
                    if (mem_test_counter < 8'hFF) begin
                        mem_test_counter <= mem_test_counter + 8'h1;
                        mem_test_addr <= mem_test_counter[9:0];
                        mem_test_data <= {24'h0, mem_test_counter};
                        
                        // Memory write/read test
                        if (mem_write_i) begin
                            // Simulate memory write
                            mem_data_o <= mem_test_data;
                        end else if (mem_read_i) begin
                            // Simulate memory read
                            mem_data_o <= mem_test_data;
                        end
                    end else begin
                        mem_test_done <= 1'b1;
                        mem_test_pass <= 1'b1;
                        mem_test_active <= 1'b0;
                    end
                end
                
                TEST_INTERFACE: begin
                    // Interface test
                    test_stage <= 8'h5;
                    test_progress_o <= 8'h80;
                    interface_active <= 1'b1;
                    loopback_ready_o <= 1'b1;
                    
                    if (interface_counter < 8'hFF) begin
                        interface_counter <= interface_counter + 8'h1;
                        interface_data <= interface_counter;
                        
                        // Loopback test
                        if (loopback_enable_i && loopback_valid_i) begin
                            loopback_data_o <= loopback_data_i;
                        end
                    end else begin
                        interface_done <= 1'b1;
                        interface_pass <= 1'b1;
                        interface_active <= 1'b0;
                    end
                end
                
                TEST_PERFORMANCE: begin
                    // Performance test
                    test_stage <= 8'h6;
                    test_progress_o <= 8'h90;
                    perf_active <= 1'b1;
                    
                    if (perf_counter < 16'hFFFF) begin
                        perf_counter <= perf_counter + 16'h1;
                        
                        // Performance benchmarking
                        if (perf_start_i) begin
                            perf_benchmark <= perf_benchmark_i;
                        end
                    end else begin
                        perf_done <= 1'b1;
                        perf_pass <= 1'b1;
                        perf_active <= 1'b0;
                        perf_result_o <= perf_counter;
                    end
                end
                
                TEST_VERIFICATION: begin
                    // Test verification
                    test_stage <= 8'h7;
                    test_progress_o <= 8'h95;
                    
                    // Verify all test results
                    if (bist_pass && scan_pass && mem_test_pass && interface_pass && perf_pass) begin
                        test_result_match <= 1'b1;
                        test_pass_count <= test_pass_count + 8'h1;
                    end else begin
                        test_result_match <= 1'b0;
                        test_error_count <= test_error_count + 8'h1;
                    end
                    
                    test_total_count <= test_total_count + 8'h1;
                    test_result_valid <= 1'b1;
                end
                
                TEST_REPORTING: begin
                    // Test reporting
                    test_stage <= 8'h8;
                    test_progress_o <= 8'h100;
                    test_done_o <= 1'b1;
                    
                    // Final test status
                    if (test_result_match) begin
                        test_pass_o <= 1'b1;
                        test_fail_o <= 1'b0;
                    end else begin
                        test_pass_o <= 1'b0;
                        test_fail_o <= 1'b1;
                    end
                    
                    // Update test status
                    test_status_o <= {test_error_count, test_pass_count};
                end
                
                TEST_ERROR: begin
                    // Test error state
                    test_stage <= 8'h9;
                    test_progress_o <= 8'h0;
                    test_fail_o <= 1'b1;
                    test_error_o <= 1'b1;
                    
                    // Reset test state
                    bist_active <= 1'b0;
                    scan_active <= 1'b0;
                    mem_test_active <= 1'b0;
                    interface_active <= 1'b0;
                    perf_active <= 1'b0;
                end
                
                default: begin
                    // No action
                end
            endcase
            
            // Test timeout handling
            if (test_active_o && test_timeout < test_timeout_limit) begin
                test_timeout <= test_timeout + 16'h1;
            end else if (test_timeout >= test_timeout_limit) begin
                test_timeout_flag <= 1'b1;
            end
        end
    end
    
    // Test data interface
    assign test_data_ready_o = (test_state == TEST_BIST || test_state == TEST_SCAN);
    
    // Memory interface
    assign mem_ready_o = (test_state == TEST_MEMORY);
    
    // Loopback interface
    assign loopback_ready_o = (test_state == TEST_INTERFACE);
    
    // Performance interface
    assign perf_done_o = (test_state == TEST_PERFORMANCE && perf_done);
    assign perf_pass_o = (test_state == TEST_PERFORMANCE && perf_pass);
    
    // Assertions for test protocol compliance
    // synthesis translate_off
    property test_state_transition;
        @(posedge PCLK_i) (test_state == TEST_IDLE) |-> ##[1:1000] (test_state != TEST_IDLE || !test_enable_i);
    endproperty
    
    property test_progress_increment;
        @(posedge PCLK_i) (test_state != TEST_IDLE) |-> ##[1:100] (test_progress_o > 8'h0);
    endproperty
    
    property test_timeout_handling;
        @(posedge PCLK_i) (test_timeout >= test_timeout_limit) |-> ##1 test_timeout_flag;
    endproperty
    
    property test_result_validation;
        @(posedge PCLK_i) (test_state == TEST_VERIFICATION) |-> ##[1:10] test_result_valid;
    endproperty
    
    property test_completion_reporting;
        @(posedge PCLK_i) (test_state == TEST_REPORTING) |-> ##[1:10] test_done_o;
    endproperty
    
    test_state_transition_check: assert property (test_state_transition)
        else $error("Test state transition violation");
    
    test_progress_increment_check: assert property (test_progress_increment)
        else $error("Test progress increment violation");
    
    test_timeout_handling_check: assert property (test_timeout_handling)
        else $error("Test timeout handling violation");
    
    test_result_validation_check: assert property (test_result_validation)
        else $error("Test result validation violation");
    
    test_completion_reporting_check: assert property (test_completion_reporting)
        else $error("Test completion reporting violation");
    // synthesis translate_on

endmodule 