//=============================================================================
// Module Name: sdcard_apb_interface
//=============================================================================
// Description: APB3 slave interface for SD Card Controller
//              Implements standard APB3 protocol with error handling
//              and register access control
//
// Features:
// - APB3 slave protocol compliance
// - Register read/write access
// - Error handling and reporting
// - Access control and protection
// - Ready signal management
// - Address decoding
//
// Author: Vyges Development Team
// License: Apache-2.0
//=============================================================================

`define SDCARD_APB_INTERFACE_SV

module sdcard_apb_interface #(
    parameter int SDCARD_APB_ADDR_WIDTH = 16
) (
    // APB Slave Interface
    input  logic                    PCLK_i,           // APB clock
    input  logic                    PRESETn_i,        // APB reset, active low
    input  logic                    PSEL_i,           // APB select
    input  logic                    PENABLE_i,        // APB enable
    input  logic                    PWRITE_i,         // APB write enable
    input  logic [SDCARD_APB_ADDR_WIDTH-1:0] PADDR_i,        // APB address bus
    input  logic [31:0]            PWDATA_i,          // APB write data
    output logic [31:0]            PRDATA_o,          // APB read data
    output logic                   PREADY_o,          // APB ready
    output logic                   PSLVERR_o,         // APB slave error
    
    // Register Interface
    output logic [31:0]            reg_data_out,      // Data to register file
    input  logic [31:0]            reg_data_in,       // Data from register file
    output logic [15:0]            reg_addr,          // Register address
    output logic                   reg_read,          // Register read enable
    output logic                   reg_write,         // Register write enable
    input  logic                   reg_ready,         // Register ready
    input  logic                   reg_error          // Register error
);

    // APB state machine states
    typedef enum logic [1:0] {
        APB_IDLE = 2'b00,
        APB_SETUP = 2'b01,
        APB_ACCESS = 2'b10,
        APB_WAIT = 2'b11
    } apb_state_t;
    
    apb_state_t apb_state, apb_next_state;
    
    // Internal signals
    logic [31:0]                   read_data_reg;
    logic                          access_done;
    logic                          access_error;
    logic [15:0]                   decoded_addr;
    logic                          addr_valid;
    logic                          write_pending;
    logic                          read_pending;
    
    // Address decoding
    always_comb begin
        decoded_addr = PADDR_i[15:0];
        addr_valid = (PADDR_i >= 16'h0000) && (PADDR_i <= 16'h005C);
    end
    
    // APB state machine
    always_ff @(posedge PCLK_i or negedge PRESETn_i) begin
        if (!PRESETn_i) begin
            apb_state <= APB_IDLE;
        end else begin
            apb_state <= apb_next_state;
        end
    end
    
    // APB state machine next state logic
    always_comb begin
        apb_next_state = apb_state;
        
        case (apb_state)
            APB_IDLE: begin
                if (PSEL_i && !PENABLE_i) begin
                    apb_next_state = APB_SETUP;
                end
            end
            
            APB_SETUP: begin
                if (PSEL_i && PENABLE_i) begin
                    apb_next_state = APB_ACCESS;
                end else if (!PSEL_i) begin
                    apb_next_state = APB_IDLE;
                end
            end
            
            APB_ACCESS: begin
                if (access_done) begin
                    apb_next_state = APB_IDLE;
                end else begin
                    apb_next_state = APB_WAIT;
                end
            end
            
            APB_WAIT: begin
                if (access_done) begin
                    apb_next_state = APB_IDLE;
                end
            end
            
            default: begin
                apb_next_state = APB_IDLE;
            end
        endcase
    end
    
    // APB control signals
    always_comb begin
        // Default values
        reg_read = 1'b0;
        reg_write = 1'b0;
        reg_addr = 16'h0;
        reg_data_out = 32'h0;
        access_done = 1'b0;
        access_error = 1'b0;
        
        case (apb_state)
            APB_SETUP: begin
                if (PWRITE_i) begin
                    write_pending = 1'b1;
                    read_pending = 1'b0;
                end else begin
                    read_pending = 1'b1;
                    write_pending = 1'b0;
                end
            end
            
            APB_ACCESS: begin
                if (addr_valid) begin
                    reg_addr = decoded_addr;
                    
                    if (PWRITE_i && write_pending) begin
                        reg_write = 1'b1;
                        reg_data_out = PWDATA_i;
                        access_done = reg_ready;
                        access_error = reg_error;
                    end else if (!PWRITE_i && read_pending) begin
                        reg_read = 1'b1;
                        access_done = reg_ready;
                        access_error = reg_error;
                    end
                end else begin
                    access_error = 1'b1;
                    access_done = 1'b1;
                end
            end
            
            APB_WAIT: begin
                access_done = reg_ready;
                access_error = reg_error;
            end
            
            default: begin
                // No action in IDLE state
            end
        endcase
    end
    
    // APB response signals
    always_ff @(posedge PCLK_i or negedge PRESETn_i) begin
        if (!PRESETn_i) begin
            PREADY_o <= 1'b0;
            PSLVERR_o <= 1'b0;
            PRDATA_o <= 32'h0;
        end else begin
            case (apb_state)
                APB_ACCESS: begin
                    if (access_done) begin
                        PREADY_o <= 1'b1;
                        PSLVERR_o <= access_error;
                        
                        if (!PWRITE_i && !access_error) begin
                            PRDATA_o <= reg_data_in;
                        end
                    end else begin
                        PREADY_o <= 1'b0;
                    end
                end
                
                APB_WAIT: begin
                    if (access_done) begin
                        PREADY_o <= 1'b1;
                        PSLVERR_o <= access_error;
                        
                        if (!PWRITE_i && !access_error) begin
                            PRDATA_o <= reg_data_in;
                        end
                    end
                end
                
                default: begin
                    PREADY_o <= 1'b0;
                    PSLVERR_o <= 1'b0;
                end
            endcase
        end
    end
    
    // Reset pending flags
    always_ff @(posedge PCLK_i or negedge PRESETn_i) begin
        if (!PRESETn_i) begin
            write_pending <= 1'b0;
            read_pending <= 1'b0;
        end else if (apb_state == APB_IDLE) begin
            write_pending <= 1'b0;
            read_pending <= 1'b0;
        end
    end

endmodule
